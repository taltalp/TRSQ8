`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date: 2017/08/17 00:56:26
// Module Name: prom
// Project Name: TRSQ8
//////////////////////////////////////////////////////////////////////////////////


module prom (
    input CLK_ip,
    input [12:0] ADDR_ip,
    output [14:0] DATA_op);

    assign DATA_op = 
        ADDR_ip==13'd0 ? 15'b010111000000000: // 
        ADDR_ip==13'd1 ? 15'b010110010000100: // 
        ADDR_ip==13'd2 ? 15'b010111011111111: // 
        ADDR_ip==13'd3 ? 15'b010110010000100: // 
        ADDR_ip==13'd4 ? 15'b110000000000000: // 
        ADDR_ip==13'd5 ? 15'b000000100000000: // 
                         15'b000000000000000;
endmodule