`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date: 2017/08/17 00:56:26
// Module Name: prom
// Project Name: TRSQ8
//////////////////////////////////////////////////////////////////////////////////


module prom (
    input CLK_ip,
    input [12:0] ADDR_ip,
    output [14:0] DATA_op);

    assign DATA_op = 
        ADDR_ip==13'd0 ? 15'b010111000000001: // 
        ADDR_ip==13'd1 ? 15'b010110000001010: // 
        ADDR_ip==13'd2 ? 15'b010111010101010: // 
        ADDR_ip==13'd3 ? 15'b010110010000010: // 
        ADDR_ip==13'd4 ? 15'b010111000010000: // 
        ADDR_ip==13'd5 ? 15'b010110010000000: // 
        ADDR_ip==13'd6 ? 15'b010110110000000: // 
        ADDR_ip==13'd7 ? 15'b010011100001010: // 
        ADDR_ip==13'd8 ? 15'b000010100000000: // 
        ADDR_ip==13'd9 ? 15'b110000000000110: // 
        ADDR_ip==13'd10 ? 15'b110000000000100: // 
        ADDR_ip==13'd11 ? 15'b000000100000000: // 
                           15'b000000000000000;
endmodule